module top(
  input wire reset,
  input wire clock
);
endmodule

